module bram_image_memory #(
    parameter int DATA_WIDTH = 8,
    parameter int ADDR_WIDTH = 10  // 2^10=1024 >= 28*28
) (
    input  logic                  clk,
    input  logic                  write_en,
    input  logic [ADDR_WIDTH-1:0] write_addr,
    input  logic [DATA_WIDTH-1:0] write_data,
    input  logic [ADDR_WIDTH-1:0] read_addr,
    output logic [DATA_WIDTH-1:0] read_data
);
    logic [DATA_WIDTH-1:0] memory [0:(1<<ADDR_WIDTH)-1];

    always_ff @(posedge clk) begin
        if (write_en) memory[write_addr] <= write_data;
        read_data <= memory[read_addr];
    end
endmodule
